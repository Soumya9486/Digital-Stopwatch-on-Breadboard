CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 0 1 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
24 C:\Program Files\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 1386 471 0 1 11
0 5
0
0 0 23408 0
2 0V
-6 -16 8 -8
4 Stop
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
45326.1 0
0
13 Logic Switch~
5 549 697 0 1 11
0 10
0
0 0 23408 0
2 0V
-6 -16 8 -8
5 Reset
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
45326.1 1
0
7 Pulser~
4 1386 409 0 10 12
0 2 84 3 85 0 0 1 1 1
8
0
0 0 6704 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3124 0 0
2
45326.1 2
0
9 2-In AND~
219 1456 461 0 3 22
0 3 5 9
0
0 0 2672 0
6 74LS08
-21 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3421 0 0
2
45326.1 3
0
8 2-In OR~
219 906 611 0 3 22
0 13 10 12
0
0 0 2672 0
6 74LS32
-21 -24 21 -16
4 U14B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8157 0 0
2
45326.1 5
0
8 2-In OR~
219 446 541 0 3 22
0 15 10 14
0
0 0 2672 0
6 74LS32
-21 -24 21 -16
4 U14A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5572 0 0
2
45326.1 6
0
9 2-In AND~
219 474 446 0 3 22
0 17 16 15
0
0 0 2672 0
6 74LS08
-21 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8901 0 0
2
45326.1 7
0
6 74LS47
187 231 255 0 14 29
0 23 22 21 20 24 24 32 33 34
35 36 37 38 24
0
0 0 6896 0
6 74LS47
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
7361 0 0
2
45326.1 8
0
6 74LS47
187 369 258 0 14 29
0 19 17 16 18 8 8 25 26 27
28 29 30 31 8
0
0 0 6896 0
6 74LS47
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
45326.1 9
0
9 CA 7-Seg~
184 386 109 0 18 19
10 38 37 36 35 34 33 32 86 11
0 0 0 0 0 0 2 2 1
0
0 0 23152 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
45326.1 10
0
9 CA 7-Seg~
184 231 109 0 18 19
10 31 30 29 28 27 26 25 87 11
0 0 0 0 0 0 2 2 1
0
0 0 23152 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3472 0 0
2
45326.1 11
0
6 74LS90
107 377 448 0 10 21
0 2 88 14 14 23 18 19 17 16
18
0
0 0 6896 0
6 74LS90
-21 -51 21 -43
2 U7
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
45326.1 12
0
6 74LS90
107 238 449 0 10 21
0 2 89 14 14 13 20 23 22 21
20
0
0 0 6896 0
6 74LS90
-21 -51 21 -43
2 U8
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
45326.1 13
0
6 74LS90
107 710 451 0 10 21
0 2 90 12 12 4 43 46 45 44
43
0
0 0 6896 0
6 74LS90
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
45326.1 14
0
6 74LS90
107 849 450 0 10 21
0 2 91 12 12 46 41 42 40 39
41
0
0 0 6896 0
6 74LS90
-21 -51 21 -43
2 U4
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3835 0 0
2
45326.1 15
0
6 74LS90
107 1088 447 0 10 21
0 2 2 10 10 9 53 50 51 52
53
0
0 0 6896 0
6 74LS90
-21 -51 21 -43
2 U5
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
45326.1 16
0
6 74LS90
107 1225 448 0 10 21
0 2 2 10 10 50 49 4 47 48
49
0
0 0 6896 0
6 74LS90
-21 -51 21 -43
2 U6
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
5616 0 0
2
45326.1 17
0
9 CA 7-Seg~
184 703 98 0 18 19
10 76 75 74 73 72 71 70 92 11
0 0 0 0 0 0 2 2 1
0
0 0 23152 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9323 0 0
2
45326.1 18
0
9 CA 7-Seg~
184 838 102 0 18 19
10 83 82 81 80 79 78 77 93 11
0 0 0 0 0 0 2 2 1
0
0 0 23152 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
317 0 0
2
45326.1 19
0
6 74LS47
187 841 260 0 14 29
0 42 40 39 41 7 7 70 71 72
73 74 75 76 7
0
0 0 6896 0
6 74LS47
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
3108 0 0
2
45326.1 20
0
6 74LS47
187 703 257 0 14 29
0 46 45 44 43 55 55 77 78 79
80 81 82 83 55
0
0 0 6896 0
6 74LS47
-21 -60 21 -52
3 U10
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
4299 0 0
2
45326.1 21
0
9 CA 7-Seg~
184 1076 101 0 18 19
10 62 61 60 59 58 57 56 94 11
0 0 0 0 2 2 0 2 1
0
0 0 23152 0
5 REDCA
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9672 0 0
2
45326.1 22
0
9 CA 7-Seg~
184 1218 102 0 18 19
10 69 68 67 66 65 64 63 95 11
0 0 0 0 0 0 2 2 1
0
0 0 23152 0
5 REDCA
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7876 0 0
2
45326.1 23
0
6 74LS47
187 1220 264 0 14 29
0 4 47 48 49 6 6 56 57 58
59 60 61 62 6
0
0 0 6896 0
6 74LS47
-21 -60 21 -52
3 U11
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
45326.1 24
0
6 74LS47
187 1082 261 0 14 29
0 50 51 52 53 54 54 63 64 65
66 67 68 69 54
0
0 0 6896 0
6 74LS47
-21 -60 21 -52
3 U12
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 0 1 0 0 0
1 U
9172 0 0
2
45326.1 25
0
8 Battery~
219 1441 116 0 2 5
0 11 2
0
0 0 2928 0
1 5
19 -2 26 6
2 V3
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
45326.1 26
0
7 Ground~
168 1442 217 0 1 3
0 2
0
0 0 55408 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
45326.1 27
0
9 2-In AND~
219 946 448 0 3 22
0 40 39 13
0
0 0 2672 0
6 74LS08
-21 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7678 0 0
2
45326.1 28
0
9 Resistor~
219 455 318 0 2 5
0 11 8
0
0 0 2928 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
45326.1 29
0
9 Resistor~
219 162 323 0 2 5
0 11 24
0
0 0 2928 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
45326.1 30
0
9 Resistor~
219 634 325 0 2 5
0 11 55
0
0 0 2928 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
45326.1 31
0
9 Resistor~
219 927 320 0 2 5
0 11 7
0
0 0 2928 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
45326.1 32
0
9 Resistor~
219 1016 321 0 2 5
0 11 54
0
0 0 2928 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
45326.1 33
0
9 Resistor~
219 1301 331 0 2 5
0 11 6
0
0 0 2928 90
2 1k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
45326.1 34
0
146
2 0 2 0 0 8192 0 17 0 0 10 4
1193 430
1183 430
1183 416
1189 416
2 0 2 0 0 0 0 16 0 0 11 4
1056 429
1046 429
1046 418
1051 418
3 1 3 0 0 8320 0 3 4 0 0 4
1410 400
1425 400
1425 452
1432 452
0 5 4 0 0 12416 0 0 14 89 0 6
1267 421
1309 421
1309 521
647 521
647 469
672 469
1 2 5 0 0 8320 0 1 4 0 0 3
1398 471
1398 470
1432 470
2 0 6 0 0 4096 0 34 0 0 106 2
1301 313
1289 313
2 0 7 0 0 8192 0 32 0 0 111 3
927 302
927 305
911 305
2 0 8 0 0 8192 0 29 0 0 49 3
455 300
455 303
443 303
0 0 2 0 0 8192 0 0 0 10 87 5
1188 395
1188 371
1406 371
1406 189
1442 189
0 1 2 0 0 0 0 0 17 11 0 4
1050 395
1189 395
1189 421
1193 421
0 1 2 0 0 4096 0 0 16 12 0 4
817 395
1051 395
1051 420
1056 420
0 1 2 0 0 0 0 0 15 13 0 3
678 395
817 395
817 423
0 1 2 0 0 4224 0 0 14 14 0 3
336 395
678 395
678 424
1 1 2 0 0 0 0 13 12 0 0 6
206 422
190 422
190 395
336 395
336 421
345 421
3 5 9 0 0 12416 0 4 16 0 0 6
1477 461
1509 461
1509 506
1035 506
1035 465
1050 465
1 2 5 0 0 0 0 1 4 0 0 3
1398 471
1398 470
1432 470
1 0 10 0 0 4096 0 2 0 0 18 4
561 697
757 697
757 646
798 646
0 0 10 0 0 12288 0 0 0 0 19 5
1215 611
1008 611
1008 653
798 653
798 617
2 2 10 0 0 12416 0 6 5 0 0 6
433 550
406 550
406 617
803 617
803 620
893 620
0 1 11 0 0 8192 0 0 26 100 0 4
1356 65
1356 48
1441 48
1441 103
0 0 10 0 0 0 0 0 0 18 86 7
1209 611
1209 606
1261 606
1261 602
1277 602
1277 553
1185 553
3 0 12 0 0 12288 0 5 0 0 26 4
939 611
955 611
955 539
808 539
1 0 13 0 0 4096 0 5 0 0 28 3
893 602
870 602
870 580
0 3 14 0 0 8192 0 0 6 27 0 5
306 547
306 634
507 634
507 541
479 541
3 1 15 0 0 12416 0 7 6 0 0 6
495 446
517 446
517 510
402 510
402 532
433 532
0 0 12 0 0 12416 0 0 0 69 70 5
663 442
629 442
629 539
808 539
808 450
0 0 14 0 0 8320 0 0 0 32 31 5
337 448
337 547
135 547
135 440
191 440
5 3 13 0 0 12416 0 13 28 0 0 5
200 467
178 467
178 580
967 580
967 448
0 9 11 0 0 8192 0 0 19 103 0 3
624 64
624 66
838 66
0 0 11 0 0 0 0 0 0 47 68 3
152 65
152 56
231 56
4 3 14 0 0 0 0 13 13 0 0 4
206 449
191 449
191 440
206 440
4 3 14 0 0 0 0 12 12 0 0 4
345 448
334 448
334 439
345 439
0 2 16 0 0 8192 0 0 7 36 0 3
428 456
428 455
450 455
0 1 17 0 0 8192 0 0 7 37 0 3
420 439
420 437
450 437
4 0 18 0 0 12416 0 9 0 0 43 6
337 249
321 249
321 359
438 359
438 475
421 475
3 9 16 0 0 8320 0 9 12 0 0 6
337 240
315 240
315 364
428 364
428 457
409 457
2 8 17 0 0 8320 0 9 12 0 0 6
337 231
311 231
311 369
420 369
420 439
409 439
1 7 19 0 0 8320 0 9 12 0 0 6
337 222
307 222
307 373
414 373
414 421
409 421
4 0 20 0 0 12416 0 8 0 0 45 6
199 246
143 246
143 380
303 380
303 476
286 476
3 9 21 0 0 8320 0 8 13 0 0 6
199 237
158 237
158 367
280 367
280 458
270 458
2 8 22 0 0 8320 0 8 13 0 0 6
199 228
176 228
176 357
288 357
288 440
270 440
1 0 23 0 0 8320 0 8 0 0 44 5
199 219
183 219
183 353
297 353
297 422
6 10 18 0 0 0 0 12 12 0 0 6
339 475
323 475
323 505
421 505
421 475
409 475
7 5 23 0 0 0 0 13 12 0 0 4
270 422
311 422
311 466
339 466
6 10 20 0 0 0 0 13 13 0 0 6
200 476
188 476
188 502
286 502
286 476
270 476
1 9 11 0 0 8192 0 29 11 0 0 5
455 336
495 336
495 58
231 58
231 73
1 0 11 0 0 8192 0 30 0 0 0 3
162 341
152 341
152 59
6 0 8 0 0 0 0 9 0 0 50 2
337 303
327 303
2 0 8 0 0 8192 0 29 0 0 50 3
455 300
455 303
412 303
5 14 8 0 0 12416 0 9 9 0 0 6
337 294
327 294
327 319
412 319
412 303
401 303
14 0 24 0 0 12416 0 8 0 0 52 5
263 300
271 300
271 312
194 312
194 300
6 0 24 0 0 0 0 8 0 0 53 3
199 300
189 300
189 291
2 5 24 0 0 0 0 30 8 0 0 3
162 305
162 291
199 291
7 7 25 0 0 8320 0 11 9 0 0 5
246 145
246 172
446 172
446 222
407 222
6 8 26 0 0 8320 0 11 9 0 0 5
240 145
240 176
441 176
441 231
407 231
5 9 27 0 0 8320 0 11 9 0 0 5
234 145
234 180
435 180
435 240
407 240
4 10 28 0 0 8320 0 11 9 0 0 5
228 145
228 184
429 184
429 249
407 249
3 11 29 0 0 8320 0 11 9 0 0 5
222 145
222 188
422 188
422 258
407 258
2 12 30 0 0 8320 0 11 9 0 0 5
216 145
216 192
417 192
417 267
407 267
1 13 31 0 0 8320 0 11 9 0 0 5
210 145
210 196
413 196
413 276
407 276
7 7 32 0 0 8320 0 10 8 0 0 5
401 145
401 158
308 158
308 219
269 219
6 8 33 0 0 8320 0 10 8 0 0 5
395 145
395 163
303 163
303 228
269 228
5 9 34 0 0 8320 0 10 8 0 0 5
389 145
389 168
296 168
296 237
269 237
4 10 35 0 0 8320 0 10 8 0 0 5
383 145
383 173
290 173
290 246
269 246
3 11 36 0 0 8320 0 10 8 0 0 5
377 145
377 177
286 177
286 255
269 255
2 12 37 0 0 8320 0 10 8 0 0 5
371 145
371 182
280 182
280 264
269 264
13 1 38 0 0 12416 0 8 10 0 0 5
269 273
275 273
275 187
365 187
365 145
9 9 11 0 0 0 0 10 11 0 0 5
386 73
231 73
231 56
231 56
231 73
4 3 12 0 0 0 0 14 14 0 0 4
678 451
663 451
663 442
678 442
4 3 12 0 0 0 0 15 15 0 0 4
817 450
805 450
805 441
817 441
0 2 39 0 0 8192 0 0 28 74 0 3
900 458
900 457
922 457
0 1 40 0 0 8192 0 0 28 75 0 3
892 441
892 439
922 439
4 0 41 0 0 12416 0 20 0 0 81 6
809 251
793 251
793 361
910 361
910 477
893 477
3 9 39 0 0 8320 0 20 15 0 0 6
809 242
787 242
787 366
900 366
900 459
881 459
2 8 40 0 0 8320 0 20 15 0 0 6
809 233
783 233
783 371
892 371
892 441
881 441
1 7 42 0 0 8320 0 20 15 0 0 6
809 224
779 224
779 375
886 375
886 423
881 423
4 0 43 0 0 12416 0 21 0 0 83 6
671 248
615 248
615 382
775 382
775 478
758 478
3 9 44 0 0 8320 0 21 14 0 0 6
671 239
630 239
630 369
752 369
752 460
742 460
2 8 45 0 0 8320 0 21 14 0 0 6
671 230
648 230
648 359
760 359
760 442
742 442
1 0 46 0 0 8320 0 21 0 0 82 5
671 221
655 221
655 355
769 355
769 424
6 10 41 0 0 0 0 15 15 0 0 6
811 477
795 477
795 507
893 507
893 477
881 477
7 5 46 0 0 0 0 14 15 0 0 4
742 424
783 424
783 468
811 468
6 10 43 0 0 0 0 14 14 0 0 6
672 478
660 478
660 504
758 504
758 478
742 478
4 0 10 0 0 0 0 16 0 0 86 3
1056 447
1042 447
1042 438
4 0 10 0 0 0 0 17 0 0 86 2
1193 448
1186 448
3 3 10 0 0 128 0 16 17 0 0 6
1056 438
1022 438
1022 553
1186 553
1186 439
1193 439
0 1 2 0 0 0 0 0 27 88 0 2
1442 179
1442 211
1 2 2 0 0 0 0 3 26 0 0 9
1362 400
1353 400
1353 375
1458 375
1458 401
1501 401
1501 179
1441 179
1441 127
1 7 4 0 0 0 0 24 17 0 0 6
1188 228
1164 228
1164 353
1267 353
1267 421
1257 421
2 8 47 0 0 8320 0 24 17 0 0 6
1188 237
1170 237
1170 345
1273 345
1273 439
1257 439
3 9 48 0 0 16512 0 24 17 0 0 6
1188 246
1179 246
1179 338
1278 338
1278 457
1257 457
4 0 49 0 0 16512 0 24 0 0 97 6
1188 255
1182 255
1182 334
1285 334
1285 476
1272 476
1 0 50 0 0 8320 0 25 0 0 98 5
1050 225
1005 225
1005 354
1123 354
1123 420
2 8 51 0 0 12416 0 25 16 0 0 6
1050 234
1010 234
1010 351
1130 351
1130 438
1120 438
3 9 52 0 0 16512 0 25 16 0 0 6
1050 243
1041 243
1041 344
1137 344
1137 456
1120 456
4 0 53 0 0 16512 0 25 0 0 99 6
1050 252
1045 252
1045 339
1143 339
1143 474
1125 474
6 10 49 0 0 0 0 17 17 0 0 6
1187 475
1175 475
1175 494
1272 494
1272 475
1257 475
7 5 50 0 0 0 0 16 17 0 0 4
1120 420
1154 420
1154 466
1187 466
6 10 53 0 0 0 0 16 16 0 0 6
1050 474
1043 474
1043 494
1125 494
1125 474
1120 474
1 9 11 0 0 8192 0 34 22 0 0 5
1301 349
1356 349
1356 64
1076 64
1076 65
1 0 11 0 0 0 0 33 0 0 145 3
1016 339
995 339
995 60
1 0 11 0 0 0 0 32 0 0 145 3
927 338
967 338
967 60
1 0 11 0 0 0 0 31 0 0 46 5
634 343
624 343
624 61
495 61
495 59
6 0 6 0 0 4096 0 24 0 0 106 2
1188 309
1174 309
14 0 6 0 0 4096 0 24 0 0 106 3
1252 309
1273 309
1273 313
5 2 6 0 0 12416 0 24 34 0 0 6
1188 300
1174 300
1174 323
1273 323
1273 313
1301 313
14 6 54 0 0 8320 0 25 25 0 0 4
1114 306
1114 322
1050 322
1050 306
5 0 54 0 0 0 0 25 0 0 109 3
1050 297
1035 297
1035 306
2 6 54 0 0 0 0 33 25 0 0 3
1016 303
1016 306
1050 306
6 0 7 0 0 0 0 20 0 0 112 2
809 305
799 305
2 0 7 0 0 8192 0 32 0 0 112 3
927 302
927 305
884 305
5 14 7 0 0 12416 0 20 20 0 0 6
809 296
799 296
799 321
884 321
884 305
873 305
14 0 55 0 0 12416 0 21 0 0 114 5
735 302
743 302
743 314
666 314
666 302
6 0 55 0 0 0 0 21 0 0 115 3
671 302
661 302
661 293
2 5 55 0 0 0 0 31 21 0 0 3
634 307
634 293
671 293
7 7 56 0 0 8320 0 22 24 0 0 5
1091 137
1091 178
1297 178
1297 228
1258 228
6 8 57 0 0 8320 0 22 24 0 0 5
1085 137
1085 182
1292 182
1292 237
1258 237
5 9 58 0 0 8320 0 22 24 0 0 5
1079 137
1079 186
1286 186
1286 246
1258 246
4 10 59 0 0 8320 0 22 24 0 0 5
1073 137
1073 190
1280 190
1280 255
1258 255
3 11 60 0 0 8320 0 22 24 0 0 5
1067 137
1067 194
1273 194
1273 264
1258 264
2 12 61 0 0 8320 0 22 24 0 0 5
1061 137
1061 198
1268 198
1268 273
1258 273
1 13 62 0 0 8320 0 22 24 0 0 5
1055 137
1055 202
1264 202
1264 282
1258 282
7 7 63 0 0 8320 0 23 25 0 0 5
1233 138
1233 164
1159 164
1159 225
1120 225
6 8 64 0 0 8320 0 23 25 0 0 5
1227 138
1227 169
1154 169
1154 234
1120 234
5 9 65 0 0 8320 0 23 25 0 0 5
1221 138
1221 174
1147 174
1147 243
1120 243
4 10 66 0 0 8320 0 23 25 0 0 5
1215 138
1215 179
1141 179
1141 252
1120 252
3 11 67 0 0 12416 0 23 25 0 0 5
1209 138
1209 183
1137 183
1137 261
1120 261
2 12 68 0 0 12416 0 23 25 0 0 5
1203 138
1203 188
1131 188
1131 270
1120 270
13 1 69 0 0 8320 0 25 23 0 0 5
1120 279
1126 279
1126 193
1197 193
1197 138
9 9 11 0 0 0 0 23 22 0 0 3
1218 66
1218 65
1076 65
7 7 70 0 0 8320 0 18 20 0 0 5
718 134
718 174
918 174
918 224
879 224
6 8 71 0 0 8320 0 18 20 0 0 5
712 134
712 178
913 178
913 233
879 233
5 9 72 0 0 8320 0 18 20 0 0 5
706 134
706 182
907 182
907 242
879 242
4 10 73 0 0 8320 0 18 20 0 0 5
700 134
700 186
901 186
901 251
879 251
3 11 74 0 0 8320 0 18 20 0 0 5
694 134
694 190
894 190
894 260
879 260
2 12 75 0 0 8320 0 18 20 0 0 5
688 134
688 194
889 194
889 269
879 269
1 13 76 0 0 8320 0 18 20 0 0 5
682 134
682 198
885 198
885 278
879 278
7 7 77 0 0 8320 0 19 21 0 0 5
853 138
853 160
780 160
780 221
741 221
6 8 78 0 0 8320 0 19 21 0 0 5
847 138
847 165
775 165
775 230
741 230
5 9 79 0 0 8320 0 19 21 0 0 5
841 138
841 170
768 170
768 239
741 239
4 10 80 0 0 8320 0 19 21 0 0 5
835 138
835 175
762 175
762 248
741 248
3 11 81 0 0 12416 0 19 21 0 0 5
829 138
829 179
758 179
758 257
741 257
2 12 82 0 0 12416 0 19 21 0 0 5
823 138
823 184
752 184
752 266
741 266
13 1 83 0 0 8320 0 21 19 0 0 5
741 275
747 275
747 189
817 189
817 138
9 9 11 0 0 8320 0 18 23 0 0 4
703 62
703 60
1218 60
1218 66
9 9 11 0 0 0 0 19 18 0 0 3
838 66
838 62
703 62
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1098 23 1199 47
1108 31 1188 47
10 Milisecond
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
738 18 807 42
748 26 796 42
6 Second
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
273 21 342 45
283 29 331 45
6 Minute
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
